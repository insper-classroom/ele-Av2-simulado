-- gray.vhd
-- Q1

Library ieee;
use ieee.std_logic_1164.all;

entity gray is
	port(
		b:      in STD_LOGIC_VECTOR(2 downto 0);
    g:      out STD_LOGIC_VECTOR(2 downto 0)
	);
end entity;

architecture rtl of gray is

begin


end architecture;
