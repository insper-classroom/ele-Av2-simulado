library IEEE; 
use IEEE.STD_LOGIC_1164.ALL;

entity fullsub is
	port ( 
			a, B, C:   in  STD_LOGIC;
			resultado, vemum:   out  STD_LOGIC);
end entity;

architecture rtl of fullsub is

begin

end;